module part4(LEDR, SW, KEY);

	input [2:0] SW;
	input [1:0] KEY;
	output [0:0] LEDR;
	
	wire 




endmodule